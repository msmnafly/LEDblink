// ********************************************************************************************************************
//
// PROJECT      :  LED Blink 
// PRODUCT      :   
// FILE         :   
// AUTHOR       :  Mohamed Nafly	
// DESCRIPTION  :  
// ********************************************************************************************************************

`timescale 1ns / 1ps

module top
#(
//---------------------------------------------------------------------------------------------------------------------
// parameter definitions
//---------------------------------------------------------------------------------------------------------------------
)(
//---------------------------------------------------------------------------------------------------------------------
// I/O signals
//---------------------------------------------------------------------------------------------------------------------
input clk,
output [1:0] LED
);

divider wrapper(
.clk(clk),
.divide(LED[0]),
.divide2(LED[1])
);
//---------------------------------------------------------------------------------------------------------------------
// Global constant headers
//---------------------------------------------------------------------------------------------------------------------

//---------------------------------------------------------------------------------------------------------------------
// localparam definitions
//---------------------------------------------------------------------------------------------------------------------

//---------------------------------------------------------------------------------------------------------------------
// Internal wires and registers
//---------------------------------------------------------------------------------------------------------------------
	
//---------------------------------------------------------------------------------------------------------------------
// Implementation
//---------------------------------------------------------------------------------------------------------------------




endmodule
