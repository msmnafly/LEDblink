// ********************************************************************************************************************
//
// PROJECT      :  LED Blink_clock divider 
// PRODUCT      :   
// FILE         :  divider.v 
// AUTHOR       :  Mohamed Nafly	
// DESCRIPTION  :   
// ********************************************************************************************************************

`timescale 1ns / 1ps

module divider
#(
//---------------------------------------------------------------------------------------------------------------------
// parameter definitions
//---------------------------------------------------------------------------------------------------------------------
)(
//---------------------------------------------------------------------------------------------------------------------
// I/O signals
//---------------------------------------------------------------------------------------------------------------------
input clk,
output reg divide = 0,
output reg divide2 = 1'b1
);

//---------------------------------------------------------------------------------------------------------------------
// Global constant headers
//---------------------------------------------------------------------------------------------------------------------
integer counter_value = 0; //32bit register
//---------------------------------------------------------------------------------------------------------------------
// localparam definitions
//---------------------------------------------------------------------------------------------------------------------
localparam div_value = 49999999;
//---------------------------------------------------------------------------------------------------------------------
// Internal wires and registers
//---------------------------------------------------------------------------------------------------------------------
	
//---------------------------------------------------------------------------------------------------------------------
// Implementation
//---------------------------------------------------------------------------------------------------------------------
always@ (posedge clk)
begin
	if (counter_value == div_value)
		counter_value <= 0;	//reset value

	else
		counter_value <= counter_value+1; //count up

end			

always@ (posedge clk)
begin
	if (counter_value == div_value)begin
		divide <= ~divide; //flip the signal 
		divide2 <= ~divide2;
	end	
	else begin
		divide <= divide; //store value	
		divide2 <= divide2;
	end	
end
endmodule
